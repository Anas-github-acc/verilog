module not_gate_xor(
    input a,
    output y
);

    xor(y, a, 1'b1);

endmodule
